module test
(
	input 	clk,
	input		reset_n,
	
	output	s
);

assign	s = 1'b0;

endmodule
