module decoder3_8 (
    input   wire            in1,
    input   wire            in2,
    input   wire            in3,
    
    output  reg     [7:0]   out
);

always @(*) begin
    case({in3,in2,in1})
        3'b000 : out = 0000_0001;
        3'b001 : out = 0000_0010;
        3'b010 : out = 0000_0100;
        3'b011 : out = 0000_1000;
        3'b100 : out = 0001_0000;
        3'b101 : out = 0010_0000;
        3'b110 : out = 0100_0000;
        3'b111 : out = 1000_0000;
        default : out = 0000_0001;
    endcase
end

endmodule