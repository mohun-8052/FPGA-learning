`timescale 1ns/1ns

module tb_mux8_1();

reg [2:0]   sel;
reg [7:0]   in;

wire        out;



endmodule